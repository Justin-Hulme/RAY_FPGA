inv_rom[1] = 16'sd32767;
inv_rom[2] = 16'sd32767;
inv_rom[3] = 16'sd32767;
inv_rom[4] = 16'sd32767;
inv_rom[5] = 16'sd32767;
inv_rom[6] = 16'sd32767;
inv_rom[7] = 16'sd32767;
inv_rom[8] = 16'sd32767;
inv_rom[9] = 16'sd32767;
inv_rom[10] = 16'sd32767;
inv_rom[11] = 16'sd32767;
inv_rom[12] = 16'sd32767;
inv_rom[13] = 16'sd32767;
inv_rom[14] = 16'sd32767;
inv_rom[15] = 16'sd32767;
inv_rom[16] = 16'sd32767;
inv_rom[17] = 16'sd32767;
inv_rom[18] = 16'sd32767;
inv_rom[19] = 16'sd32767;
inv_rom[20] = 16'sd32767;
inv_rom[21] = 16'sd32767;
inv_rom[22] = 16'sd32767;
inv_rom[23] = 16'sd32767;
inv_rom[24] = 16'sd32767;
inv_rom[25] = 16'sd32767;
inv_rom[26] = 16'sd32767;
inv_rom[27] = 16'sd32767;
inv_rom[28] = 16'sd32767;
inv_rom[29] = 16'sd32767;
inv_rom[30] = 16'sd32767;
inv_rom[31] = 16'sd32767;
inv_rom[32] = 16'sd32767;
inv_rom[33] = 16'sd32767;
inv_rom[34] = 16'sd32767;
inv_rom[35] = 16'sd32767;
inv_rom[36] = 16'sd32767;
inv_rom[37] = 16'sd32767;
inv_rom[38] = 16'sd32767;
inv_rom[39] = 16'sd32767;
inv_rom[40] = 16'sd32767;
inv_rom[41] = 16'sd32767;
inv_rom[42] = 16'sd32767;
inv_rom[43] = 16'sd32767;
inv_rom[44] = 16'sd32767;
inv_rom[45] = 16'sd32767;
inv_rom[46] = 16'sd32767;
inv_rom[47] = 16'sd32767;
inv_rom[48] = 16'sd32767;
inv_rom[49] = 16'sd32767;
inv_rom[50] = 16'sd32767;
inv_rom[51] = 16'sd32767;
inv_rom[52] = 16'sd32767;
inv_rom[53] = 16'sd32767;
inv_rom[54] = 16'sd32767;
inv_rom[55] = 16'sd32767;
inv_rom[56] = 16'sd32767;
inv_rom[57] = 16'sd32767;
inv_rom[58] = 16'sd32767;
inv_rom[59] = 16'sd32767;
inv_rom[60] = 16'sd32767;
inv_rom[61] = 16'sd32767;
inv_rom[62] = 16'sd32767;
inv_rom[63] = 16'sd32767;
inv_rom[64] = 16'sd32767;
inv_rom[65] = 16'sd32767;
inv_rom[66] = 16'sd32767;
inv_rom[67] = 16'sd32767;
inv_rom[68] = 16'sd32767;
inv_rom[69] = 16'sd32767;
inv_rom[70] = 16'sd32767;
inv_rom[71] = 16'sd32767;
inv_rom[72] = 16'sd32767;
inv_rom[73] = 16'sd32767;
inv_rom[74] = 16'sd32767;
inv_rom[75] = 16'sd32767;
inv_rom[76] = 16'sd32767;
inv_rom[77] = 16'sd32767;
inv_rom[78] = 16'sd32767;
inv_rom[79] = 16'sd32767;
inv_rom[80] = 16'sd32767;
inv_rom[81] = 16'sd32767;
inv_rom[82] = 16'sd32767;
inv_rom[83] = 16'sd32767;
inv_rom[84] = 16'sd32767;
inv_rom[85] = 16'sd32767;
inv_rom[86] = 16'sd32767;
inv_rom[87] = 16'sd32767;
inv_rom[88] = 16'sd32767;
inv_rom[89] = 16'sd32767;
inv_rom[90] = 16'sd32767;
inv_rom[91] = 16'sd32767;
inv_rom[92] = 16'sd32767;
inv_rom[93] = 16'sd32767;
inv_rom[94] = 16'sd32767;
inv_rom[95] = 16'sd32767;
inv_rom[96] = 16'sd32767;
inv_rom[97] = 16'sd32767;
inv_rom[98] = 16'sd32767;
inv_rom[99] = 16'sd32767;
inv_rom[100] = 16'sd32767;
inv_rom[101] = 16'sd32767;
inv_rom[102] = 16'sd32767;
inv_rom[103] = 16'sd32767;
inv_rom[104] = 16'sd32767;
inv_rom[105] = 16'sd32767;
inv_rom[106] = 16'sd32767;
inv_rom[107] = 16'sd32767;
inv_rom[108] = 16'sd32767;
inv_rom[109] = 16'sd32767;
inv_rom[110] = 16'sd32767;
inv_rom[111] = 16'sd32767;
inv_rom[112] = 16'sd32767;
inv_rom[113] = 16'sd32767;
inv_rom[114] = 16'sd32767;
inv_rom[115] = 16'sd32767;
inv_rom[116] = 16'sd32767;
inv_rom[117] = 16'sd32767;
inv_rom[118] = 16'sd32767;
inv_rom[119] = 16'sd32767;
inv_rom[120] = 16'sd32767;
inv_rom[121] = 16'sd32767;
inv_rom[122] = 16'sd32767;
inv_rom[123] = 16'sd32767;
inv_rom[124] = 16'sd32767;
inv_rom[125] = 16'sd32767;
inv_rom[126] = 16'sd32767;
inv_rom[127] = 16'sd32767;
inv_rom[128] = 16'sd32767;
inv_rom[129] = 16'sd32514;
inv_rom[130] = 16'sd32264;
inv_rom[131] = 16'sd32018;
inv_rom[132] = 16'sd31775;
inv_rom[133] = 16'sd31536;
inv_rom[134] = 16'sd31301;
inv_rom[135] = 16'sd31069;
inv_rom[136] = 16'sd30840;
inv_rom[137] = 16'sd30615;
inv_rom[138] = 16'sd30394;
inv_rom[139] = 16'sd30175;
inv_rom[140] = 16'sd29959;
inv_rom[141] = 16'sd29747;
inv_rom[142] = 16'sd29537;
inv_rom[143] = 16'sd29331;
inv_rom[144] = 16'sd29127;
inv_rom[145] = 16'sd28926;
inv_rom[146] = 16'sd28728;
inv_rom[147] = 16'sd28533;
inv_rom[148] = 16'sd28340;
inv_rom[149] = 16'sd28150;
inv_rom[150] = 16'sd27962;
inv_rom[151] = 16'sd27777;
inv_rom[152] = 16'sd27594;
inv_rom[153] = 16'sd27414;
inv_rom[154] = 16'sd27236;
inv_rom[155] = 16'sd27060;
inv_rom[156] = 16'sd26887;
inv_rom[157] = 16'sd26715;
inv_rom[158] = 16'sd26546;
inv_rom[159] = 16'sd26379;
inv_rom[160] = 16'sd26214;
inv_rom[161] = 16'sd26052;
inv_rom[162] = 16'sd25891;
inv_rom[163] = 16'sd25732;
inv_rom[164] = 16'sd25575;
inv_rom[165] = 16'sd25420;
inv_rom[166] = 16'sd25267;
inv_rom[167] = 16'sd25116;
inv_rom[168] = 16'sd24966;
inv_rom[169] = 16'sd24818;
inv_rom[170] = 16'sd24672;
inv_rom[171] = 16'sd24528;
inv_rom[172] = 16'sd24385;
inv_rom[173] = 16'sd24245;
inv_rom[174] = 16'sd24105;
inv_rom[175] = 16'sd23967;
inv_rom[176] = 16'sd23831;
inv_rom[177] = 16'sd23697;
inv_rom[178] = 16'sd23564;
inv_rom[179] = 16'sd23432;
inv_rom[180] = 16'sd23302;
inv_rom[181] = 16'sd23173;
inv_rom[182] = 16'sd23046;
inv_rom[183] = 16'sd22920;
inv_rom[184] = 16'sd22795;
inv_rom[185] = 16'sd22672;
inv_rom[186] = 16'sd22550;
inv_rom[187] = 16'sd22429;
inv_rom[188] = 16'sd22310;
inv_rom[189] = 16'sd22192;
inv_rom[190] = 16'sd22075;
inv_rom[191] = 16'sd21960;
inv_rom[192] = 16'sd21845;
inv_rom[193] = 16'sd21732;
inv_rom[194] = 16'sd21620;
inv_rom[195] = 16'sd21509;
inv_rom[196] = 16'sd21400;
inv_rom[197] = 16'sd21291;
inv_rom[198] = 16'sd21183;
inv_rom[199] = 16'sd21077;
inv_rom[200] = 16'sd20972;
inv_rom[201] = 16'sd20867;
inv_rom[202] = 16'sd20764;
inv_rom[203] = 16'sd20662;
inv_rom[204] = 16'sd20560;
inv_rom[205] = 16'sd20460;
inv_rom[206] = 16'sd20361;
inv_rom[207] = 16'sd20262;
inv_rom[208] = 16'sd20165;
inv_rom[209] = 16'sd20068;
inv_rom[210] = 16'sd19973;
inv_rom[211] = 16'sd19878;
inv_rom[212] = 16'sd19784;
inv_rom[213] = 16'sd19692;
inv_rom[214] = 16'sd19600;
inv_rom[215] = 16'sd19508;
inv_rom[216] = 16'sd19418;
inv_rom[217] = 16'sd19329;
inv_rom[218] = 16'sd19240;
inv_rom[219] = 16'sd19152;
inv_rom[220] = 16'sd19065;
inv_rom[221] = 16'sd18979;
inv_rom[222] = 16'sd18893;
inv_rom[223] = 16'sd18809;
inv_rom[224] = 16'sd18725;
inv_rom[225] = 16'sd18641;
inv_rom[226] = 16'sd18559;
inv_rom[227] = 16'sd18477;
inv_rom[228] = 16'sd18396;
inv_rom[229] = 16'sd18316;
inv_rom[230] = 16'sd18236;
inv_rom[231] = 16'sd18157;
inv_rom[232] = 16'sd18079;
inv_rom[233] = 16'sd18001;
inv_rom[234] = 16'sd17924;
inv_rom[235] = 16'sd17848;
inv_rom[236] = 16'sd17772;
inv_rom[237] = 16'sd17697;
inv_rom[238] = 16'sd17623;
inv_rom[239] = 16'sd17549;
inv_rom[240] = 16'sd17476;
inv_rom[241] = 16'sd17404;
inv_rom[242] = 16'sd17332;
inv_rom[243] = 16'sd17261;
inv_rom[244] = 16'sd17190;
inv_rom[245] = 16'sd17120;
inv_rom[246] = 16'sd17050;
inv_rom[247] = 16'sd16981;
inv_rom[248] = 16'sd16913;
inv_rom[249] = 16'sd16845;
inv_rom[250] = 16'sd16777;
inv_rom[251] = 16'sd16710;
inv_rom[252] = 16'sd16644;
inv_rom[253] = 16'sd16578;
inv_rom[254] = 16'sd16513;
inv_rom[255] = 16'sd16448;
inv_rom[0] = 16'sd32767;

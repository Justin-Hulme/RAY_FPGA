sin_rom[0] = 16'sd0;
sin_rom[1] = 16'sd402;
sin_rom[2] = 16'sd804;
sin_rom[3] = 16'sd1205;
sin_rom[4] = 16'sd1606;
sin_rom[5] = 16'sd2006;
sin_rom[6] = 16'sd2404;
sin_rom[7] = 16'sd2801;
sin_rom[8] = 16'sd3196;
sin_rom[9] = 16'sd3590;
sin_rom[10] = 16'sd3981;
sin_rom[11] = 16'sd4370;
sin_rom[12] = 16'sd4756;
sin_rom[13] = 16'sd5139;
sin_rom[14] = 16'sd5520;
sin_rom[15] = 16'sd5897;
sin_rom[16] = 16'sd6270;
sin_rom[17] = 16'sd6639;
sin_rom[18] = 16'sd7005;
sin_rom[19] = 16'sd7366;
sin_rom[20] = 16'sd7723;
sin_rom[21] = 16'sd8076;
sin_rom[22] = 16'sd8423;
sin_rom[23] = 16'sd8765;
sin_rom[24] = 16'sd9102;
sin_rom[25] = 16'sd9434;
sin_rom[26] = 16'sd9760;
sin_rom[27] = 16'sd10080;
sin_rom[28] = 16'sd10394;
sin_rom[29] = 16'sd10702;
sin_rom[30] = 16'sd11003;
sin_rom[31] = 16'sd11297;
sin_rom[32] = 16'sd11585;
sin_rom[33] = 16'sd11866;
sin_rom[34] = 16'sd12140;
sin_rom[35] = 16'sd12406;
sin_rom[36] = 16'sd12665;
sin_rom[37] = 16'sd12916;
sin_rom[38] = 16'sd13160;
sin_rom[39] = 16'sd13395;
sin_rom[40] = 16'sd13623;
sin_rom[41] = 16'sd13842;
sin_rom[42] = 16'sd14053;
sin_rom[43] = 16'sd14256;
sin_rom[44] = 16'sd14449;
sin_rom[45] = 16'sd14635;
sin_rom[46] = 16'sd14811;
sin_rom[47] = 16'sd14978;
sin_rom[48] = 16'sd15137;
sin_rom[49] = 16'sd15286;
sin_rom[50] = 16'sd15426;
sin_rom[51] = 16'sd15557;
sin_rom[52] = 16'sd15679;
sin_rom[53] = 16'sd15791;
sin_rom[54] = 16'sd15893;
sin_rom[55] = 16'sd15986;
sin_rom[56] = 16'sd16069;
sin_rom[57] = 16'sd16143;
sin_rom[58] = 16'sd16207;
sin_rom[59] = 16'sd16261;
sin_rom[60] = 16'sd16305;
sin_rom[61] = 16'sd16340;
sin_rom[62] = 16'sd16364;
sin_rom[63] = 16'sd16379;
sin_rom[64] = 16'sd16384;
sin_rom[65] = 16'sd16379;
sin_rom[66] = 16'sd16364;
sin_rom[67] = 16'sd16340;
sin_rom[68] = 16'sd16305;
sin_rom[69] = 16'sd16261;
sin_rom[70] = 16'sd16207;
sin_rom[71] = 16'sd16143;
sin_rom[72] = 16'sd16069;
sin_rom[73] = 16'sd15986;
sin_rom[74] = 16'sd15893;
sin_rom[75] = 16'sd15791;
sin_rom[76] = 16'sd15679;
sin_rom[77] = 16'sd15557;
sin_rom[78] = 16'sd15426;
sin_rom[79] = 16'sd15286;
sin_rom[80] = 16'sd15137;
sin_rom[81] = 16'sd14978;
sin_rom[82] = 16'sd14811;
sin_rom[83] = 16'sd14635;
sin_rom[84] = 16'sd14449;
sin_rom[85] = 16'sd14256;
sin_rom[86] = 16'sd14053;
sin_rom[87] = 16'sd13842;
sin_rom[88] = 16'sd13623;
sin_rom[89] = 16'sd13395;
sin_rom[90] = 16'sd13160;
sin_rom[91] = 16'sd12916;
sin_rom[92] = 16'sd12665;
sin_rom[93] = 16'sd12406;
sin_rom[94] = 16'sd12140;
sin_rom[95] = 16'sd11866;
sin_rom[96] = 16'sd11585;
sin_rom[97] = 16'sd11297;
sin_rom[98] = 16'sd11003;
sin_rom[99] = 16'sd10702;
sin_rom[100] = 16'sd10394;
sin_rom[101] = 16'sd10080;
sin_rom[102] = 16'sd9760;
sin_rom[103] = 16'sd9434;
sin_rom[104] = 16'sd9102;
sin_rom[105] = 16'sd8765;
sin_rom[106] = 16'sd8423;
sin_rom[107] = 16'sd8076;
sin_rom[108] = 16'sd7723;
sin_rom[109] = 16'sd7366;
sin_rom[110] = 16'sd7005;
sin_rom[111] = 16'sd6639;
sin_rom[112] = 16'sd6270;
sin_rom[113] = 16'sd5897;
sin_rom[114] = 16'sd5520;
sin_rom[115] = 16'sd5139;
sin_rom[116] = 16'sd4756;
sin_rom[117] = 16'sd4370;
sin_rom[118] = 16'sd3981;
sin_rom[119] = 16'sd3590;
sin_rom[120] = 16'sd3196;
sin_rom[121] = 16'sd2801;
sin_rom[122] = 16'sd2404;
sin_rom[123] = 16'sd2006;
sin_rom[124] = 16'sd1606;
sin_rom[125] = 16'sd1205;
sin_rom[126] = 16'sd804;
sin_rom[127] = 16'sd402;
sin_rom[128] = 16'sd0;
sin_rom[129] = -16'sd402;
sin_rom[130] = -16'sd804;
sin_rom[131] = -16'sd1205;
sin_rom[132] = -16'sd1606;
sin_rom[133] = -16'sd2006;
sin_rom[134] = -16'sd2404;
sin_rom[135] = -16'sd2801;
sin_rom[136] = -16'sd3196;
sin_rom[137] = -16'sd3590;
sin_rom[138] = -16'sd3981;
sin_rom[139] = -16'sd4370;
sin_rom[140] = -16'sd4756;
sin_rom[141] = -16'sd5139;
sin_rom[142] = -16'sd5520;
sin_rom[143] = -16'sd5897;
sin_rom[144] = -16'sd6270;
sin_rom[145] = -16'sd6639;
sin_rom[146] = -16'sd7005;
sin_rom[147] = -16'sd7366;
sin_rom[148] = -16'sd7723;
sin_rom[149] = -16'sd8076;
sin_rom[150] = -16'sd8423;
sin_rom[151] = -16'sd8765;
sin_rom[152] = -16'sd9102;
sin_rom[153] = -16'sd9434;
sin_rom[154] = -16'sd9760;
sin_rom[155] = -16'sd10080;
sin_rom[156] = -16'sd10394;
sin_rom[157] = -16'sd10702;
sin_rom[158] = -16'sd11003;
sin_rom[159] = -16'sd11297;
sin_rom[160] = -16'sd11585;
sin_rom[161] = -16'sd11866;
sin_rom[162] = -16'sd12140;
sin_rom[163] = -16'sd12406;
sin_rom[164] = -16'sd12665;
sin_rom[165] = -16'sd12916;
sin_rom[166] = -16'sd13160;
sin_rom[167] = -16'sd13395;
sin_rom[168] = -16'sd13623;
sin_rom[169] = -16'sd13842;
sin_rom[170] = -16'sd14053;
sin_rom[171] = -16'sd14256;
sin_rom[172] = -16'sd14449;
sin_rom[173] = -16'sd14635;
sin_rom[174] = -16'sd14811;
sin_rom[175] = -16'sd14978;
sin_rom[176] = -16'sd15137;
sin_rom[177] = -16'sd15286;
sin_rom[178] = -16'sd15426;
sin_rom[179] = -16'sd15557;
sin_rom[180] = -16'sd15679;
sin_rom[181] = -16'sd15791;
sin_rom[182] = -16'sd15893;
sin_rom[183] = -16'sd15986;
sin_rom[184] = -16'sd16069;
sin_rom[185] = -16'sd16143;
sin_rom[186] = -16'sd16207;
sin_rom[187] = -16'sd16261;
sin_rom[188] = -16'sd16305;
sin_rom[189] = -16'sd16340;
sin_rom[190] = -16'sd16364;
sin_rom[191] = -16'sd16379;
sin_rom[192] = -16'sd16384;
sin_rom[193] = -16'sd16379;
sin_rom[194] = -16'sd16364;
sin_rom[195] = -16'sd16340;
sin_rom[196] = -16'sd16305;
sin_rom[197] = -16'sd16261;
sin_rom[198] = -16'sd16207;
sin_rom[199] = -16'sd16143;
sin_rom[200] = -16'sd16069;
sin_rom[201] = -16'sd15986;
sin_rom[202] = -16'sd15893;
sin_rom[203] = -16'sd15791;
sin_rom[204] = -16'sd15679;
sin_rom[205] = -16'sd15557;
sin_rom[206] = -16'sd15426;
sin_rom[207] = -16'sd15286;
sin_rom[208] = -16'sd15137;
sin_rom[209] = -16'sd14978;
sin_rom[210] = -16'sd14811;
sin_rom[211] = -16'sd14635;
sin_rom[212] = -16'sd14449;
sin_rom[213] = -16'sd14256;
sin_rom[214] = -16'sd14053;
sin_rom[215] = -16'sd13842;
sin_rom[216] = -16'sd13623;
sin_rom[217] = -16'sd13395;
sin_rom[218] = -16'sd13160;
sin_rom[219] = -16'sd12916;
sin_rom[220] = -16'sd12665;
sin_rom[221] = -16'sd12406;
sin_rom[222] = -16'sd12140;
sin_rom[223] = -16'sd11866;
sin_rom[224] = -16'sd11585;
sin_rom[225] = -16'sd11297;
sin_rom[226] = -16'sd11003;
sin_rom[227] = -16'sd10702;
sin_rom[228] = -16'sd10394;
sin_rom[229] = -16'sd10080;
sin_rom[230] = -16'sd9760;
sin_rom[231] = -16'sd9434;
sin_rom[232] = -16'sd9102;
sin_rom[233] = -16'sd8765;
sin_rom[234] = -16'sd8423;
sin_rom[235] = -16'sd8076;
sin_rom[236] = -16'sd7723;
sin_rom[237] = -16'sd7366;
sin_rom[238] = -16'sd7005;
sin_rom[239] = -16'sd6639;
sin_rom[240] = -16'sd6270;
sin_rom[241] = -16'sd5897;
sin_rom[242] = -16'sd5520;
sin_rom[243] = -16'sd5139;
sin_rom[244] = -16'sd4756;
sin_rom[245] = -16'sd4370;
sin_rom[246] = -16'sd3981;
sin_rom[247] = -16'sd3590;
sin_rom[248] = -16'sd3196;
sin_rom[249] = -16'sd2801;
sin_rom[250] = -16'sd2404;
sin_rom[251] = -16'sd2006;
sin_rom[252] = -16'sd1606;
sin_rom[253] = -16'sd1205;
sin_rom[254] = -16'sd804;
sin_rom[255] = -16'sd402;
